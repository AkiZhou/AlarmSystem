library ieee;
	use ieee.std_logic_1164.all;
	
entity DispFrac is
	port (HEX0, HEX1, HEX2, HEX3 : out std_logic_vector(6 downto 0));
end DispFrac;